module dec2to4(W,en, Y);
/*
endmodule
*/